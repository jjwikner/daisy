.include /sw/cadence/libraries/cmos065_522/IO65LPHVT_SF_2V5_50A_7M4X0Y2Z_7.0/physical/IO65LPHVT_SF_2V5_50A_7M4X0Y2Z.cdl
